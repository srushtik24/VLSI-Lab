magic
tech scmos
timestamp 1642154095
<< nwell >>
rect -8 7 18 23
<< polysilicon >>
rect -3 13 1 15
rect 9 13 13 15
rect -3 -3 1 9
rect 9 -3 13 9
rect -1 -7 1 -3
rect 11 -7 13 -3
rect -3 -10 1 -7
rect 9 -10 13 -7
rect -3 -16 1 -14
rect 9 -16 13 -14
<< ndiffusion >>
rect -4 -14 -3 -10
rect 1 -14 9 -10
rect 13 -14 14 -10
<< pdiffusion >>
rect -4 9 -3 13
rect 1 9 3 13
rect 7 9 9 13
rect 13 9 14 13
<< metal1 >>
rect -12 21 18 22
rect -12 17 3 21
rect 7 17 18 21
rect -8 13 -4 17
rect 14 13 18 17
rect 3 5 7 9
rect 3 1 22 5
rect -9 -7 -5 -3
rect 3 -7 7 -3
rect 14 -10 18 1
rect -8 -18 -4 -14
rect -12 -22 -8 -18
<< ntransistor >>
rect -3 -14 1 -10
rect 9 -14 13 -10
<< ptransistor >>
rect -3 9 1 13
rect 9 9 13 13
<< polycontact >>
rect -5 -7 -1 -3
rect 7 -7 11 -3
<< ndcontact >>
rect -8 -14 -4 -10
rect 14 -14 18 -10
<< pdcontact >>
rect -8 9 -4 13
rect 3 9 7 13
rect 14 9 18 13
<< psubstratepcontact >>
rect -8 -22 -4 -18
<< nsubstratencontact >>
rect 3 17 7 21
<< labels >>
rlabel metal1 -11 20 -11 20 4 vdd
rlabel metal1 -11 -19 -11 -19 2 gnd
rlabel metal1 -9 -7 -9 -3 3 A
rlabel metal1 3 -7 3 -3 1 B
rlabel metal1 22 1 22 5 7 Out
<< end >>
